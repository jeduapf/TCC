* C:\Users\jedua\Desktop\UNICAMP\UNICAMP_2022\2sem2022\TCC\Pspice_Python\Circuits\Circuito5_cargas_RLC.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 13 18:18:53 2022



** Analysis setup **
.tran 1us 150ms 0 1us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Circuito5_cargas_RLC.net"
.INC "Circuito5_cargas_RLC.als"


.probe/CSDF N($N_0029) 
.probe/CSDF I(R_Rcorrente) 


.END
