* C:\Users\jedua\Desktop\UNICAMP\UNICAMP_2022\2sem2022\TCC\Pspice_Python\Circuits\Circuito4_cargar_diferentes.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 13 18:18:23 2022



** Analysis setup **
.tran 1us 150ms 0 1us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Circuito4_cargar_diferentes.net"
.INC "Circuito4_cargar_diferentes.als"


.probe/CSDF N(A) 
.probe/CSDF I(R_Rcorrente) 


.END
